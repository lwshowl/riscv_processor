module icache #(way)(
);


// each cache line is 64 bytes long
// for a set associative cache , each way is 4k bytes large
ram #(WIDTH=8,ENTRY=4028)()



endmodule