module dcache (
    ports
);
    
endmodule