module axi_ctl(
    input r_req1,
    input [63:0] r_addr1,
    output r_data1;
    output r_ready;

    input r_req2,
    input r_addr2,
    output r_data2,

    input w_req1,
    input w_addr1,
    input w_data1,
);


endmodule